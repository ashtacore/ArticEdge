`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: Jay Runyan
// 
// Create Date: 07/20/2024 09:15:48 PM
// Design Name: ArcticEdge
// Module Name: top
// Project Name: arctic_edge_core
// Target Devices: Nexys A7-100T
// Tool Versions: Vivado 2024.1
// Description: Building my own RISC-V core in System Verilog
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module cpu_core(
    input wire clk,                   // Board clock
);

endmodule